// niosiisystem.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module niosiisystem (
		output wire        adc_sclk,      //       adc.sclk
		output wire        adc_cs_n,      //          .cs_n
		input  wire        adc_dout,      //          .dout
		output wire        adc_din,       //          .din
		input  wire        clk_clk,       //       clk.clk
		output wire [15:0] gpio_export,   //      gpio.export
		output wire [9:0]  ledr_export,   //      ledr.export
		input  wire        reset_reset,   //     reset.reset
		output wire [12:0] sdram_addr,    //     sdram.addr
		output wire [1:0]  sdram_ba,      //          .ba
		output wire        sdram_cas_n,   //          .cas_n
		output wire        sdram_cke,     //          .cke
		output wire        sdram_cs_n,    //          .cs_n
		inout  wire [15:0] sdram_dq,      //          .dq
		output wire [1:0]  sdram_dqm,     //          .dqm
		output wire        sdram_ras_n,   //          .ras_n
		output wire        sdram_we_n,    //          .we_n
		output wire        sdram_clk_clk, // sdram_clk.clk
		input  wire [9:0]  switch_export  //    switch.export
	);

	wire         sys_sdram_pll_0_sys_clk_clk;                                 // sys_sdram_pll_0:sys_clk_clk -> [DRAM:clk, GPIO:clk, IMEM:clk, LEDR:clk, SW:clk, adc_0:clock, irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:sys_sdram_pll_0_sys_clk_clk, nios2_gen2_0:clk, rst_controller:clk, rst_controller_001:clk, sysid_qsys_0:clock, timer_0:clk, timer_1:clk]
	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [26:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [26:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire  [31:0] mm_interconnect_0_adc_0_adc_slave_readdata;                  // adc_0:readdata -> mm_interconnect_0:adc_0_adc_slave_readdata
	wire         mm_interconnect_0_adc_0_adc_slave_waitrequest;               // adc_0:waitrequest -> mm_interconnect_0:adc_0_adc_slave_waitrequest
	wire   [2:0] mm_interconnect_0_adc_0_adc_slave_address;                   // mm_interconnect_0:adc_0_adc_slave_address -> adc_0:address
	wire         mm_interconnect_0_adc_0_adc_slave_read;                      // mm_interconnect_0:adc_0_adc_slave_read -> adc_0:read
	wire         mm_interconnect_0_adc_0_adc_slave_write;                     // mm_interconnect_0:adc_0_adc_slave_write -> adc_0:write
	wire  [31:0] mm_interconnect_0_adc_0_adc_slave_writedata;                 // mm_interconnect_0:adc_0_adc_slave_writedata -> adc_0:writedata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;       // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;        // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_imem_s1_chipselect;                        // mm_interconnect_0:IMEM_s1_chipselect -> IMEM:chipselect
	wire  [31:0] mm_interconnect_0_imem_s1_readdata;                          // IMEM:readdata -> mm_interconnect_0:IMEM_s1_readdata
	wire  [15:0] mm_interconnect_0_imem_s1_address;                           // mm_interconnect_0:IMEM_s1_address -> IMEM:address
	wire   [3:0] mm_interconnect_0_imem_s1_byteenable;                        // mm_interconnect_0:IMEM_s1_byteenable -> IMEM:byteenable
	wire         mm_interconnect_0_imem_s1_write;                             // mm_interconnect_0:IMEM_s1_write -> IMEM:write
	wire  [31:0] mm_interconnect_0_imem_s1_writedata;                         // mm_interconnect_0:IMEM_s1_writedata -> IMEM:writedata
	wire         mm_interconnect_0_imem_s1_clken;                             // mm_interconnect_0:IMEM_s1_clken -> IMEM:clken
	wire         mm_interconnect_0_dram_s1_chipselect;                        // mm_interconnect_0:DRAM_s1_chipselect -> DRAM:az_cs
	wire  [15:0] mm_interconnect_0_dram_s1_readdata;                          // DRAM:za_data -> mm_interconnect_0:DRAM_s1_readdata
	wire         mm_interconnect_0_dram_s1_waitrequest;                       // DRAM:za_waitrequest -> mm_interconnect_0:DRAM_s1_waitrequest
	wire  [24:0] mm_interconnect_0_dram_s1_address;                           // mm_interconnect_0:DRAM_s1_address -> DRAM:az_addr
	wire         mm_interconnect_0_dram_s1_read;                              // mm_interconnect_0:DRAM_s1_read -> DRAM:az_rd_n
	wire   [1:0] mm_interconnect_0_dram_s1_byteenable;                        // mm_interconnect_0:DRAM_s1_byteenable -> DRAM:az_be_n
	wire         mm_interconnect_0_dram_s1_readdatavalid;                     // DRAM:za_valid -> mm_interconnect_0:DRAM_s1_readdatavalid
	wire         mm_interconnect_0_dram_s1_write;                             // mm_interconnect_0:DRAM_s1_write -> DRAM:az_wr_n
	wire  [15:0] mm_interconnect_0_dram_s1_writedata;                         // mm_interconnect_0:DRAM_s1_writedata -> DRAM:az_data
	wire  [31:0] mm_interconnect_0_sw_s1_readdata;                            // SW:readdata -> mm_interconnect_0:SW_s1_readdata
	wire   [1:0] mm_interconnect_0_sw_s1_address;                             // mm_interconnect_0:SW_s1_address -> SW:address
	wire         mm_interconnect_0_ledr_s1_chipselect;                        // mm_interconnect_0:LEDR_s1_chipselect -> LEDR:chipselect
	wire  [31:0] mm_interconnect_0_ledr_s1_readdata;                          // LEDR:readdata -> mm_interconnect_0:LEDR_s1_readdata
	wire   [1:0] mm_interconnect_0_ledr_s1_address;                           // mm_interconnect_0:LEDR_s1_address -> LEDR:address
	wire         mm_interconnect_0_ledr_s1_write;                             // mm_interconnect_0:LEDR_s1_write -> LEDR:write_n
	wire  [31:0] mm_interconnect_0_ledr_s1_writedata;                         // mm_interconnect_0:LEDR_s1_writedata -> LEDR:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                     // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                        // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                          // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                      // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_timer_1_s1_chipselect;                     // mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	wire  [15:0] mm_interconnect_0_timer_1_s1_readdata;                       // timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_1_s1_address;                        // mm_interconnect_0:timer_1_s1_address -> timer_1:address
	wire         mm_interconnect_0_timer_1_s1_write;                          // mm_interconnect_0:timer_1_s1_write -> timer_1:write_n
	wire  [15:0] mm_interconnect_0_timer_1_s1_writedata;                      // mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	wire         mm_interconnect_0_gpio_s1_chipselect;                        // mm_interconnect_0:GPIO_s1_chipselect -> GPIO:chipselect
	wire  [31:0] mm_interconnect_0_gpio_s1_readdata;                          // GPIO:readdata -> mm_interconnect_0:GPIO_s1_readdata
	wire   [1:0] mm_interconnect_0_gpio_s1_address;                           // mm_interconnect_0:GPIO_s1_address -> GPIO:address
	wire         mm_interconnect_0_gpio_s1_write;                             // mm_interconnect_0:GPIO_s1_write -> GPIO:write_n
	wire  [31:0] mm_interconnect_0_gpio_s1_writedata;                         // mm_interconnect_0:GPIO_s1_writedata -> GPIO:writedata
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // timer_1:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // timer_0:irq -> irq_mapper:receiver2_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [DRAM:reset_n, GPIO:reset_n, IMEM:reset, LEDR:reset_n, SW:reset_n, adc_0:reset, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, rst_translator:in_reset, sysid_qsys_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [IMEM:reset_req, nios2_gen2_0:reset_req, rst_translator:reset_req_in]
	wire         sys_sdram_pll_0_reset_source_reset;                          // sys_sdram_pll_0:reset_source_reset -> [rst_controller:reset_in0, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [mm_interconnect_0:timer_0_reset_reset_bridge_in_reset_reset, timer_0:reset_n, timer_1:reset_n]
	wire         nios2_gen2_0_debug_reset_request_reset;                      // nios2_gen2_0:debug_reset_request -> rst_controller_001:reset_in0

	niosiisystem_DRAM dram (
		.clk            (sys_sdram_pll_0_sys_clk_clk),             //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),         // reset.reset_n
		.az_addr        (mm_interconnect_0_dram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_dram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_dram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_dram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_dram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_dram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_dram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_dram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_dram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                              //  wire.export
		.zs_ba          (sdram_ba),                                //      .export
		.zs_cas_n       (sdram_cas_n),                             //      .export
		.zs_cke         (sdram_cke),                               //      .export
		.zs_cs_n        (sdram_cs_n),                              //      .export
		.zs_dq          (sdram_dq),                                //      .export
		.zs_dqm         (sdram_dqm),                               //      .export
		.zs_ras_n       (sdram_ras_n),                             //      .export
		.zs_we_n        (sdram_we_n)                               //      .export
	);

	niosiisystem_GPIO gpio (
		.clk        (sys_sdram_pll_0_sys_clk_clk),          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_gpio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gpio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gpio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gpio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gpio_s1_readdata),   //                    .readdata
		.out_port   (gpio_export)                           // external_connection.export
	);

	niosiisystem_IMEM imem (
		.clk        (sys_sdram_pll_0_sys_clk_clk),          //   clk1.clk
		.address    (mm_interconnect_0_imem_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_imem_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_imem_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_imem_s1_write),      //       .write
		.readdata   (mm_interconnect_0_imem_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_imem_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_imem_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),   //       .reset_req
		.freeze     (1'b0)                                  // (terminated)
	);

	niosiisystem_LEDR ledr (
		.clk        (sys_sdram_pll_0_sys_clk_clk),          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledr_s1_readdata),   //                    .readdata
		.out_port   (ledr_export)                           // external_connection.export
	);

	niosiisystem_SW sw (
		.clk      (sys_sdram_pll_0_sys_clk_clk),      //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_0_sw_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sw_s1_readdata), //                    .readdata
		.in_port  (switch_export)                     // external_connection.export
	);

	niosiisystem_adc_0 #(
		.board          ("DE10-Standard"),
		.board_rev      ("Autodetect"),
		.tsclk          (4),
		.numch          (7),
		.max10pllmultby (1),
		.max10plldivby  (1)
	) adc_0 (
		.clock       (sys_sdram_pll_0_sys_clk_clk),                   //                clk.clk
		.reset       (rst_controller_reset_out_reset),                //              reset.reset
		.write       (mm_interconnect_0_adc_0_adc_slave_write),       //          adc_slave.write
		.readdata    (mm_interconnect_0_adc_0_adc_slave_readdata),    //                   .readdata
		.writedata   (mm_interconnect_0_adc_0_adc_slave_writedata),   //                   .writedata
		.address     (mm_interconnect_0_adc_0_adc_slave_address),     //                   .address
		.waitrequest (mm_interconnect_0_adc_0_adc_slave_waitrequest), //                   .waitrequest
		.read        (mm_interconnect_0_adc_0_adc_slave_read),        //                   .read
		.adc_sclk    (adc_sclk),                                      // external_interface.export
		.adc_cs_n    (adc_cs_n),                                      //                   .export
		.adc_dout    (adc_dout),                                      //                   .export
		.adc_din     (adc_din)                                        //                   .export
	);

	niosiisystem_jtag_uart_0 jtag_uart_0 (
		.clk            (sys_sdram_pll_0_sys_clk_clk),                                 //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	niosiisystem_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (sys_sdram_pll_0_sys_clk_clk),                                //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	niosiisystem_sys_sdram_pll_0 sys_sdram_pll_0 (
		.ref_clk_clk        (clk_clk),                            //      ref_clk.clk
		.ref_reset_reset    (reset_reset),                        //    ref_reset.reset
		.sys_clk_clk        (sys_sdram_pll_0_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                      //    sdram_clk.clk
		.reset_source_reset (sys_sdram_pll_0_reset_source_reset)  // reset_source.reset
	);

	niosiisystem_sysid_qsys_0 sysid_qsys_0 (
		.clock    (sys_sdram_pll_0_sys_clk_clk),                           //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	niosiisystem_timer_0 timer_0 (
		.clk        (sys_sdram_pll_0_sys_clk_clk),             //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                 //   irq.irq
	);

	niosiisystem_timer_0 timer_1 (
		.clk        (sys_sdram_pll_0_sys_clk_clk),             //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	niosiisystem_mm_interconnect_0 mm_interconnect_0 (
		.sys_sdram_pll_0_sys_clk_clk                    (sys_sdram_pll_0_sys_clk_clk),                                 //                  sys_sdram_pll_0_sys_clk.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.timer_0_reset_reset_bridge_in_reset_reset      (rst_controller_001_reset_out_reset),                          //      timer_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                            //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                         //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                               //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                           //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                              //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                          //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                     //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                        //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                    //                                         .readdata
		.adc_0_adc_slave_address                        (mm_interconnect_0_adc_0_adc_slave_address),                   //                          adc_0_adc_slave.address
		.adc_0_adc_slave_write                          (mm_interconnect_0_adc_0_adc_slave_write),                     //                                         .write
		.adc_0_adc_slave_read                           (mm_interconnect_0_adc_0_adc_slave_read),                      //                                         .read
		.adc_0_adc_slave_readdata                       (mm_interconnect_0_adc_0_adc_slave_readdata),                  //                                         .readdata
		.adc_0_adc_slave_writedata                      (mm_interconnect_0_adc_0_adc_slave_writedata),                 //                                         .writedata
		.adc_0_adc_slave_waitrequest                    (mm_interconnect_0_adc_0_adc_slave_waitrequest),               //                                         .waitrequest
		.DRAM_s1_address                                (mm_interconnect_0_dram_s1_address),                           //                                  DRAM_s1.address
		.DRAM_s1_write                                  (mm_interconnect_0_dram_s1_write),                             //                                         .write
		.DRAM_s1_read                                   (mm_interconnect_0_dram_s1_read),                              //                                         .read
		.DRAM_s1_readdata                               (mm_interconnect_0_dram_s1_readdata),                          //                                         .readdata
		.DRAM_s1_writedata                              (mm_interconnect_0_dram_s1_writedata),                         //                                         .writedata
		.DRAM_s1_byteenable                             (mm_interconnect_0_dram_s1_byteenable),                        //                                         .byteenable
		.DRAM_s1_readdatavalid                          (mm_interconnect_0_dram_s1_readdatavalid),                     //                                         .readdatavalid
		.DRAM_s1_waitrequest                            (mm_interconnect_0_dram_s1_waitrequest),                       //                                         .waitrequest
		.DRAM_s1_chipselect                             (mm_interconnect_0_dram_s1_chipselect),                        //                                         .chipselect
		.GPIO_s1_address                                (mm_interconnect_0_gpio_s1_address),                           //                                  GPIO_s1.address
		.GPIO_s1_write                                  (mm_interconnect_0_gpio_s1_write),                             //                                         .write
		.GPIO_s1_readdata                               (mm_interconnect_0_gpio_s1_readdata),                          //                                         .readdata
		.GPIO_s1_writedata                              (mm_interconnect_0_gpio_s1_writedata),                         //                                         .writedata
		.GPIO_s1_chipselect                             (mm_interconnect_0_gpio_s1_chipselect),                        //                                         .chipselect
		.IMEM_s1_address                                (mm_interconnect_0_imem_s1_address),                           //                                  IMEM_s1.address
		.IMEM_s1_write                                  (mm_interconnect_0_imem_s1_write),                             //                                         .write
		.IMEM_s1_readdata                               (mm_interconnect_0_imem_s1_readdata),                          //                                         .readdata
		.IMEM_s1_writedata                              (mm_interconnect_0_imem_s1_writedata),                         //                                         .writedata
		.IMEM_s1_byteenable                             (mm_interconnect_0_imem_s1_byteenable),                        //                                         .byteenable
		.IMEM_s1_chipselect                             (mm_interconnect_0_imem_s1_chipselect),                        //                                         .chipselect
		.IMEM_s1_clken                                  (mm_interconnect_0_imem_s1_clken),                             //                                         .clken
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.LEDR_s1_address                                (mm_interconnect_0_ledr_s1_address),                           //                                  LEDR_s1.address
		.LEDR_s1_write                                  (mm_interconnect_0_ledr_s1_write),                             //                                         .write
		.LEDR_s1_readdata                               (mm_interconnect_0_ledr_s1_readdata),                          //                                         .readdata
		.LEDR_s1_writedata                              (mm_interconnect_0_ledr_s1_writedata),                         //                                         .writedata
		.LEDR_s1_chipselect                             (mm_interconnect_0_ledr_s1_chipselect),                        //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.SW_s1_address                                  (mm_interconnect_0_sw_s1_address),                             //                                    SW_s1.address
		.SW_s1_readdata                                 (mm_interconnect_0_sw_s1_readdata),                            //                                         .readdata
		.sysid_qsys_0_control_slave_address             (mm_interconnect_0_sysid_qsys_0_control_slave_address),        //               sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata            (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),       //                                         .readdata
		.timer_0_s1_address                             (mm_interconnect_0_timer_0_s1_address),                        //                               timer_0_s1.address
		.timer_0_s1_write                               (mm_interconnect_0_timer_0_s1_write),                          //                                         .write
		.timer_0_s1_readdata                            (mm_interconnect_0_timer_0_s1_readdata),                       //                                         .readdata
		.timer_0_s1_writedata                           (mm_interconnect_0_timer_0_s1_writedata),                      //                                         .writedata
		.timer_0_s1_chipselect                          (mm_interconnect_0_timer_0_s1_chipselect),                     //                                         .chipselect
		.timer_1_s1_address                             (mm_interconnect_0_timer_1_s1_address),                        //                               timer_1_s1.address
		.timer_1_s1_write                               (mm_interconnect_0_timer_1_s1_write),                          //                                         .write
		.timer_1_s1_readdata                            (mm_interconnect_0_timer_1_s1_readdata),                       //                                         .readdata
		.timer_1_s1_writedata                           (mm_interconnect_0_timer_1_s1_writedata),                      //                                         .writedata
		.timer_1_s1_chipselect                          (mm_interconnect_0_timer_1_s1_chipselect)                      //                                         .chipselect
	);

	niosiisystem_irq_mapper irq_mapper (
		.clk           (sys_sdram_pll_0_sys_clk_clk),    //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (sys_sdram_pll_0_reset_source_reset), // reset_in0.reset
		.clk            (sys_sdram_pll_0_sys_clk_clk),        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (nios2_gen2_0_debug_reset_request_reset), // reset_in0.reset
		.reset_in1      (sys_sdram_pll_0_reset_source_reset),     // reset_in1.reset
		.clk            (sys_sdram_pll_0_sys_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
